module top();
input a,b;
output reg s,c;
always(*)begin
s=a+b;
c=ab;
end
endmodule